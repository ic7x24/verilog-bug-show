`define NUM_1 8'b0101_1111;
`define NUM_2 8'h01
`define NUM_3 32'd1000000
`define NUM_3 {4'h0, 4{1'b1}}
`define NUM_5 {4'h1, 4{1'b1}}

